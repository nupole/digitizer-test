library ieee;
use ieee.std_logic_1164.all;

package types_pkg is
    type array_std_logic_vector is array(natural range<>) of std_logic_vector;
end package;
