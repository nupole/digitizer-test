library ieee;
use ieee.std_logic_1164.all;

library work;
use work.types_pkg.all;

package local_bus_interface_pkg is
    alias registers is array_std_logic_vector;
end package;
